module conv_test;


